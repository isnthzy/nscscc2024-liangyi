module DiffBridge(
    input        clock,
    input [ 7:0] coreid,
    input [ 7:0] index_0,
    input        Instrvalid_0,
    input [63:0] the_pc_0,
    input [31:0] instr_0,
    input        skip_0,
    input        is_TLBFILL_0,
    input [ 4:0] TLBFILL_index_0,
    input        is_CNTinst_0,
    input [63:0] timer_64_value_0,
    input        wen_0,
    input [ 7:0] wdest_0,
    input [63:0] wdata_0,
    input        csr_rstat_0,
    input [31:0] csr_data_0,

    input [ 7:0] index_1,
    input        Instrvalid_1,
    input [63:0] the_pc_1,
    input [31:0] instr_1,
    input        skip_1,
    input        is_TLBFILL_1,
    input [ 4:0] TLBFILL_index_1,
    input        is_CNTinst_1,
    input [63:0] timer_64_value_1,
    input        wen_1,
    input [ 7:0] wdest_1,
    input [63:0] wdata_1,
    input        csr_rstat_1,
    input [31:0] csr_data_1,

    input        excp_valid,
    input        eret,
    input [31:0] intrNo,
    input [31:0] cause,
    input [63:0] exceptionPC,
    input [31:0] exceptionInst,

    input [ 7:0] storeIndex_0,
    input [ 7:0] storeValid_0,
    input [63:0] storePaddr_0,
    input [63:0] storeVaddr_0,
    input [63:0] storeData_0,

    input [ 7:0] storeIndex_1,
    input [ 7:0] storeValid_1,
    input [63:0] storePaddr_1,
    input [63:0] storeVaddr_1,
    input [63:0] storeData_1,

    input [ 7:0] loadIndex_0,
    input [ 7:0] loadValid_0,
    input [63:0] loadPaddr_0,
    input [63:0] loadVaddr_0,

    input [ 7:0] loadIndex_1,
    input [ 7:0] loadValid_1,
    input [63:0] loadPaddr_1,
    input [63:0] loadVaddr_1,


    input [63:0] crmd,
    input [63:0] prmd,
    input [63:0] euen,
    input [63:0] ecfg,
    input [63:0] estat,
    input [63:0] era,
    input [63:0] badv,
    input [63:0] eentry,
    input [63:0] tlbidx,
    input [63:0] tlbehi,
    input [63:0] tlbelo0,
    input [63:0] tlbelo1,
    input [63:0] asid,
    input [63:0] pgdl,
    input [63:0] pgdh,
    input [63:0] save0,
    input [63:0] save1,
    input [63:0] save2,
    input [63:0] save3,
    input [63:0] tid,
    input [63:0] tcfg,
    input [63:0] tval,
    input [63:0] ticlr,
    input [63:0] llbctl,
    input [63:0] tlbrentry,
    input [63:0] dmw0,
    input [63:0] dmw1,

    input [63:0] REG_0,
    input [63:0] REG_1,
    input [63:0] REG_2,
    input [63:0] REG_3,
    input [63:0] REG_4,
    input [63:0] REG_5,
    input [63:0] REG_6,
    input [63:0] REG_7,
    input [63:0] REG_8,
    input [63:0] REG_9,
    input [63:0] REG_10,
    input [63:0] REG_11,
    input [63:0] REG_12,
    input [63:0] REG_13,
    input [63:0] REG_14,
    input [63:0] REG_15,
    input [63:0] REG_16,
    input [63:0] REG_17,
    input [63:0] REG_18,
    input [63:0] REG_19,
    input [63:0] REG_20,
    input [63:0] REG_21,
    input [63:0] REG_22,
    input [63:0] REG_23,
    input [63:0] REG_24,
    input [63:0] REG_25,
    input [63:0] REG_26,
    input [63:0] REG_27,
    input [63:0] REG_28,
    input [63:0] REG_29,
    input [63:0] REG_30,
    input [63:0] REG_31

);

DifftestInstrCommit DifftestInstrCommit_0(
    .clock              (clock          ),
    .coreid             (coreid         ),
    .index              (index_0        ),
    .valid              (Instrvalid_0   ),
    .pc                 (the_pc_0       ),
    .instr              (instr_0        ),
    .skip               (skip_0         ),
    .is_TLBFILL         (is_TLBFILL_0   ),
    .TLBFILL_index      (TLBFILL_index_0),
    .is_CNTinst         (is_CNTinst_0   ),
    .timer_64_value     (timer_64_value_0),
    .wen                (wen_0          ),
    .wdest              (wdest_0        ),
    .wdata              (wdata_0        ),
    .csr_rstat          (csr_rstat_0    ),
    .csr_data           (csr_data_0     )
);

DifftestStoreEvent DifftestStoreEvent_0(
    .clock              (clock          ),
    .coreid             (0              ),
    .index              (storeIndex_0   ),
    .valid              (storeValid_0   ),
    .storePAddr         (storePaddr_0   ),
    .storeVAddr         (storeVaddr_0   ),
    .storeData          (storeData_0    )
);

DifftestLoadEvent DifftestLoadEvent_0(
    .clock              (clock          ),
    .coreid             (0              ),
    .index              (loadIndex_0    ),
    .valid              (loadValid_0    ),
    .paddr              (loadPaddr_0    ),
    .vaddr              (loadVaddr_0    )
);

DifftestInstrCommit DifftestInstrCommit_1(
    .clock              (clock          ),
    .coreid             (coreid         ),
    .index              (index_1        ),
    .valid              (Instrvalid_1   ),
    .pc                 (the_pc_1       ),
    .instr              (instr_1        ),
    .skip               (skip_1         ),
    .is_TLBFILL         (is_TLBFILL_1   ),
    .TLBFILL_index      (TLBFILL_index_1),
    .is_CNTinst         (is_CNTinst_1   ),
    .timer_64_value     (timer_64_value_1),
    .wen                (wen_1          ),
    .wdest              (wdest_1        ),
    .wdata              (wdata_1        ),
    .csr_rstat          (csr_rstat_1    ),
    .csr_data           (csr_data_1     )
);

DifftestStoreEvent DifftestStoreEvent_1(
    .clock              (clock          ),
    .coreid             (0              ),
    .index              (storeIndex_1   ),
    .valid              (storeValid_1   ),
    .storePAddr         (storePaddr_1   ),
    .storeVAddr         (storeVaddr_1   ),
    .storeData          (storeData_1    )
);

DifftestLoadEvent DifftestLoadEvent(
    .clock              (clock          ),
    .coreid             (0              ),
    .index              (loadIndex_1    ),
    .valid              (loadValid_1    ),
    .paddr              (loadPaddr_1    ),
    .vaddr              (loadVaddr_1    )
);


DifftestExcpEvent DifftestExcpEvent(
    .clock              (clock          ),
    .coreid             (coreid         ),
    .excp_valid         (excp_valid     ),
    .eret               (eret           ),
    .intrNo             (intrNo[12:2]   ),
    .cause              (cause          ),
    .exceptionPC        (exceptionPC    ),
    .exceptionInst      (exceptionInst  )
);

DifftestTrapEvent DifftestTrapEvent(
    .clock              (clock          ),
    .coreid             (0              ),
    .valid              (0              ),
    .code               (0              ),
    .pc                 (0              ),
    .cycleCnt           (0              ),
    .instrCnt           (0              )
);

DifftestCSRRegState DifftestCSRRegState(
    .clock              (clock              ),
    .coreid             (0                  ),
    .crmd               (crmd               ),
    .prmd               (prmd               ),
    .euen               (euen               ),
    .ecfg               (ecfg               ),
    .estat              (estat              ),
    .era                (era                ),
    .badv               (badv               ),
    .eentry             (eentry             ),
    .tlbidx             (tlbidx             ),
    .tlbehi             (tlbehi             ),
    .tlbelo0            (tlbelo0            ),
    .tlbelo1            (tlbelo1            ),
    .asid               (asid               ),
    .pgdl               (pgdl               ),
    .pgdh               (pgdh               ),
    .save0              (save0              ),
    .save1              (save1              ),
    .save2              (save2              ),
    .save3              (save3              ),
    .tid                (tid                ),
    .tcfg               (tcfg               ),
    .tval               (tval               ),
    .ticlr              (ticlr              ),
    .llbctl             (llbctl             ),
    .tlbrentry          (tlbrentry          ),
    .dmw0               (dmw0               ),
    .dmw1               (dmw1               )
);

DifftestGRegState DifftestGRegState(
    .clock              (clock     ),
    .coreid             (0         ),
    .gpr_0              (0         ),
    .gpr_1              (REG_1     ),
    .gpr_2              (REG_2     ),
    .gpr_3              (REG_3     ),
    .gpr_4              (REG_4     ),
    .gpr_5              (REG_5     ),
    .gpr_6              (REG_6     ),
    .gpr_7              (REG_7     ),
    .gpr_8              (REG_8     ),
    .gpr_9              (REG_9     ),
    .gpr_10             (REG_10    ),
    .gpr_11             (REG_11    ),
    .gpr_12             (REG_12    ),
    .gpr_13             (REG_13    ),
    .gpr_14             (REG_14    ),
    .gpr_15             (REG_15    ),
    .gpr_16             (REG_16    ),
    .gpr_17             (REG_17    ),
    .gpr_18             (REG_18    ),
    .gpr_19             (REG_19    ),
    .gpr_20             (REG_20    ),
    .gpr_21             (REG_21    ),
    .gpr_22             (REG_22    ),
    .gpr_23             (REG_23    ),
    .gpr_24             (REG_24    ),
    .gpr_25             (REG_25    ),
    .gpr_26             (REG_26    ),
    .gpr_27             (REG_27    ),
    .gpr_28             (REG_28    ),
    .gpr_29             (REG_29    ),
    .gpr_30             (REG_30    ),
    .gpr_31             (REG_31    )
);

endmodule